
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h068b5899;
    ram_cell[       1] = 32'h0;  // 32'hb078a2d2;
    ram_cell[       2] = 32'h0;  // 32'hf0d2f875;
    ram_cell[       3] = 32'h0;  // 32'h45b8f052;
    ram_cell[       4] = 32'h0;  // 32'hf27c7987;
    ram_cell[       5] = 32'h0;  // 32'h74430d0b;
    ram_cell[       6] = 32'h0;  // 32'he1739a30;
    ram_cell[       7] = 32'h0;  // 32'h9b8c4edc;
    ram_cell[       8] = 32'h0;  // 32'hee8873f1;
    ram_cell[       9] = 32'h0;  // 32'hc49045fa;
    ram_cell[      10] = 32'h0;  // 32'h7cf9ed4d;
    ram_cell[      11] = 32'h0;  // 32'hc0126625;
    ram_cell[      12] = 32'h0;  // 32'h4aa649e1;
    ram_cell[      13] = 32'h0;  // 32'h0161e4b2;
    ram_cell[      14] = 32'h0;  // 32'hfbbf9b9e;
    ram_cell[      15] = 32'h0;  // 32'h3759b2f8;
    ram_cell[      16] = 32'h0;  // 32'hdfdcf7ed;
    ram_cell[      17] = 32'h0;  // 32'h36794929;
    ram_cell[      18] = 32'h0;  // 32'hc7961eb6;
    ram_cell[      19] = 32'h0;  // 32'h35f5f318;
    ram_cell[      20] = 32'h0;  // 32'hc729c403;
    ram_cell[      21] = 32'h0;  // 32'h71da519c;
    ram_cell[      22] = 32'h0;  // 32'h03261e4d;
    ram_cell[      23] = 32'h0;  // 32'h5226ed56;
    ram_cell[      24] = 32'h0;  // 32'he7aefeb1;
    ram_cell[      25] = 32'h0;  // 32'hb0a07591;
    ram_cell[      26] = 32'h0;  // 32'hff9f7bb7;
    ram_cell[      27] = 32'h0;  // 32'hf1856304;
    ram_cell[      28] = 32'h0;  // 32'he1ea00c8;
    ram_cell[      29] = 32'h0;  // 32'h833492eb;
    ram_cell[      30] = 32'h0;  // 32'hb1ec6195;
    ram_cell[      31] = 32'h0;  // 32'h8ef36c58;
    ram_cell[      32] = 32'h0;  // 32'he7a7aadc;
    ram_cell[      33] = 32'h0;  // 32'hafb3b3a9;
    ram_cell[      34] = 32'h0;  // 32'h6f017dd4;
    ram_cell[      35] = 32'h0;  // 32'hf5e90d57;
    ram_cell[      36] = 32'h0;  // 32'h43f86973;
    ram_cell[      37] = 32'h0;  // 32'h9b5b987d;
    ram_cell[      38] = 32'h0;  // 32'h92ab8200;
    ram_cell[      39] = 32'h0;  // 32'h0ef89dfb;
    ram_cell[      40] = 32'h0;  // 32'hece72196;
    ram_cell[      41] = 32'h0;  // 32'haf0fd9d0;
    ram_cell[      42] = 32'h0;  // 32'h117ebb5a;
    ram_cell[      43] = 32'h0;  // 32'h5abc0a9b;
    ram_cell[      44] = 32'h0;  // 32'he03214e7;
    ram_cell[      45] = 32'h0;  // 32'he75aa48d;
    ram_cell[      46] = 32'h0;  // 32'h37b29b81;
    ram_cell[      47] = 32'h0;  // 32'h0ada687e;
    ram_cell[      48] = 32'h0;  // 32'hb4dd5020;
    ram_cell[      49] = 32'h0;  // 32'hc70146e7;
    ram_cell[      50] = 32'h0;  // 32'h765b99bf;
    ram_cell[      51] = 32'h0;  // 32'h96c26201;
    ram_cell[      52] = 32'h0;  // 32'h86425e90;
    ram_cell[      53] = 32'h0;  // 32'h5b6864ad;
    ram_cell[      54] = 32'h0;  // 32'h7243cf6c;
    ram_cell[      55] = 32'h0;  // 32'h68bc7364;
    ram_cell[      56] = 32'h0;  // 32'ha32af3bc;
    ram_cell[      57] = 32'h0;  // 32'hb55046f5;
    ram_cell[      58] = 32'h0;  // 32'h862506db;
    ram_cell[      59] = 32'h0;  // 32'h3ebe6e97;
    ram_cell[      60] = 32'h0;  // 32'hdd331041;
    ram_cell[      61] = 32'h0;  // 32'hcc6b9ca7;
    ram_cell[      62] = 32'h0;  // 32'h73083d34;
    ram_cell[      63] = 32'h0;  // 32'hdca49c37;
    ram_cell[      64] = 32'h0;  // 32'hdcc69f49;
    ram_cell[      65] = 32'h0;  // 32'h170a64dd;
    ram_cell[      66] = 32'h0;  // 32'ha95aa2e8;
    ram_cell[      67] = 32'h0;  // 32'h21a27d3f;
    ram_cell[      68] = 32'h0;  // 32'hb9bea659;
    ram_cell[      69] = 32'h0;  // 32'h874fe083;
    ram_cell[      70] = 32'h0;  // 32'hc50dc22a;
    ram_cell[      71] = 32'h0;  // 32'h5703433e;
    ram_cell[      72] = 32'h0;  // 32'h5d5e13e9;
    ram_cell[      73] = 32'h0;  // 32'h09b16863;
    ram_cell[      74] = 32'h0;  // 32'h54ecc769;
    ram_cell[      75] = 32'h0;  // 32'h602fea69;
    ram_cell[      76] = 32'h0;  // 32'hf9dd3ecf;
    ram_cell[      77] = 32'h0;  // 32'he11926a9;
    ram_cell[      78] = 32'h0;  // 32'h2fb4a9ac;
    ram_cell[      79] = 32'h0;  // 32'h86a6fe26;
    ram_cell[      80] = 32'h0;  // 32'h19ebf52b;
    ram_cell[      81] = 32'h0;  // 32'h6a63bb3f;
    ram_cell[      82] = 32'h0;  // 32'hd2f67454;
    ram_cell[      83] = 32'h0;  // 32'habfbcef9;
    ram_cell[      84] = 32'h0;  // 32'hb082f03b;
    ram_cell[      85] = 32'h0;  // 32'h05f40a66;
    ram_cell[      86] = 32'h0;  // 32'h2c19cb69;
    ram_cell[      87] = 32'h0;  // 32'h96c432c8;
    ram_cell[      88] = 32'h0;  // 32'h5db5b1b5;
    ram_cell[      89] = 32'h0;  // 32'h44cc9de2;
    ram_cell[      90] = 32'h0;  // 32'h6399bb2d;
    ram_cell[      91] = 32'h0;  // 32'hb3f9d118;
    ram_cell[      92] = 32'h0;  // 32'h715c3a65;
    ram_cell[      93] = 32'h0;  // 32'hf6a1465d;
    ram_cell[      94] = 32'h0;  // 32'h9c516e08;
    ram_cell[      95] = 32'h0;  // 32'h50daebeb;
    ram_cell[      96] = 32'h0;  // 32'h245bf71f;
    ram_cell[      97] = 32'h0;  // 32'h1c697678;
    ram_cell[      98] = 32'h0;  // 32'ha80da9d2;
    ram_cell[      99] = 32'h0;  // 32'h12c2ae5c;
    ram_cell[     100] = 32'h0;  // 32'h90afd6c9;
    ram_cell[     101] = 32'h0;  // 32'h71939e2a;
    ram_cell[     102] = 32'h0;  // 32'h127777ba;
    ram_cell[     103] = 32'h0;  // 32'h6ab40dfd;
    ram_cell[     104] = 32'h0;  // 32'he21b19bf;
    ram_cell[     105] = 32'h0;  // 32'h61d4632f;
    ram_cell[     106] = 32'h0;  // 32'hf0af2335;
    ram_cell[     107] = 32'h0;  // 32'h1c31245a;
    ram_cell[     108] = 32'h0;  // 32'h5deb1a4c;
    ram_cell[     109] = 32'h0;  // 32'h9607c9de;
    ram_cell[     110] = 32'h0;  // 32'he5d68caf;
    ram_cell[     111] = 32'h0;  // 32'h44c964d2;
    ram_cell[     112] = 32'h0;  // 32'h8bac054c;
    ram_cell[     113] = 32'h0;  // 32'h57af0ebe;
    ram_cell[     114] = 32'h0;  // 32'h0a5770bd;
    ram_cell[     115] = 32'h0;  // 32'h22600e89;
    ram_cell[     116] = 32'h0;  // 32'h69383738;
    ram_cell[     117] = 32'h0;  // 32'he4444ae1;
    ram_cell[     118] = 32'h0;  // 32'h7e00d294;
    ram_cell[     119] = 32'h0;  // 32'h74ff3d84;
    ram_cell[     120] = 32'h0;  // 32'hc3784fbb;
    ram_cell[     121] = 32'h0;  // 32'h0c345452;
    ram_cell[     122] = 32'h0;  // 32'ha9ea3f31;
    ram_cell[     123] = 32'h0;  // 32'h2dedccbb;
    ram_cell[     124] = 32'h0;  // 32'hb13b7c80;
    ram_cell[     125] = 32'h0;  // 32'hd7d80112;
    ram_cell[     126] = 32'h0;  // 32'h96d2f984;
    ram_cell[     127] = 32'h0;  // 32'hfb789f7c;
    ram_cell[     128] = 32'h0;  // 32'hf95725fc;
    ram_cell[     129] = 32'h0;  // 32'hf6eb72c9;
    ram_cell[     130] = 32'h0;  // 32'hf990713e;
    ram_cell[     131] = 32'h0;  // 32'hd23dbde7;
    ram_cell[     132] = 32'h0;  // 32'ha2d9f5e6;
    ram_cell[     133] = 32'h0;  // 32'hd1aca98b;
    ram_cell[     134] = 32'h0;  // 32'h7d04ce45;
    ram_cell[     135] = 32'h0;  // 32'h51aab161;
    ram_cell[     136] = 32'h0;  // 32'h6062aea1;
    ram_cell[     137] = 32'h0;  // 32'h72d0cdfd;
    ram_cell[     138] = 32'h0;  // 32'h9f9573a8;
    ram_cell[     139] = 32'h0;  // 32'hc216631d;
    ram_cell[     140] = 32'h0;  // 32'hcc8189b1;
    ram_cell[     141] = 32'h0;  // 32'h4cc08f2e;
    ram_cell[     142] = 32'h0;  // 32'h122c64fa;
    ram_cell[     143] = 32'h0;  // 32'hac6889d1;
    ram_cell[     144] = 32'h0;  // 32'hb9446ea3;
    ram_cell[     145] = 32'h0;  // 32'h693efec6;
    ram_cell[     146] = 32'h0;  // 32'ha5706a6b;
    ram_cell[     147] = 32'h0;  // 32'h2afb185a;
    ram_cell[     148] = 32'h0;  // 32'h73693897;
    ram_cell[     149] = 32'h0;  // 32'hd3d0d530;
    ram_cell[     150] = 32'h0;  // 32'h52946664;
    ram_cell[     151] = 32'h0;  // 32'he9847c79;
    ram_cell[     152] = 32'h0;  // 32'hdfaa50f9;
    ram_cell[     153] = 32'h0;  // 32'hc3e8d3d1;
    ram_cell[     154] = 32'h0;  // 32'h5bb38013;
    ram_cell[     155] = 32'h0;  // 32'he78cfddd;
    ram_cell[     156] = 32'h0;  // 32'h97b04758;
    ram_cell[     157] = 32'h0;  // 32'haf8ec882;
    ram_cell[     158] = 32'h0;  // 32'h05cccb1e;
    ram_cell[     159] = 32'h0;  // 32'h49448848;
    ram_cell[     160] = 32'h0;  // 32'h23881b51;
    ram_cell[     161] = 32'h0;  // 32'hdbcda82b;
    ram_cell[     162] = 32'h0;  // 32'h989f14f1;
    ram_cell[     163] = 32'h0;  // 32'h056608c1;
    ram_cell[     164] = 32'h0;  // 32'h59b3e212;
    ram_cell[     165] = 32'h0;  // 32'h6d5d7485;
    ram_cell[     166] = 32'h0;  // 32'ha398f766;
    ram_cell[     167] = 32'h0;  // 32'h16a69884;
    ram_cell[     168] = 32'h0;  // 32'ha91bcd93;
    ram_cell[     169] = 32'h0;  // 32'h33699241;
    ram_cell[     170] = 32'h0;  // 32'h5939413f;
    ram_cell[     171] = 32'h0;  // 32'he3f71b8a;
    ram_cell[     172] = 32'h0;  // 32'h8b52d3ee;
    ram_cell[     173] = 32'h0;  // 32'h8779473f;
    ram_cell[     174] = 32'h0;  // 32'h710875cf;
    ram_cell[     175] = 32'h0;  // 32'h03ba084e;
    ram_cell[     176] = 32'h0;  // 32'h8eaf2edd;
    ram_cell[     177] = 32'h0;  // 32'h44d265c7;
    ram_cell[     178] = 32'h0;  // 32'h6ac8bbfd;
    ram_cell[     179] = 32'h0;  // 32'hd1b53c82;
    ram_cell[     180] = 32'h0;  // 32'hee9ddc52;
    ram_cell[     181] = 32'h0;  // 32'hfb362a51;
    ram_cell[     182] = 32'h0;  // 32'heade6fa3;
    ram_cell[     183] = 32'h0;  // 32'hdf1b9cf3;
    ram_cell[     184] = 32'h0;  // 32'hbf5b0993;
    ram_cell[     185] = 32'h0;  // 32'h9e492512;
    ram_cell[     186] = 32'h0;  // 32'h735b51ff;
    ram_cell[     187] = 32'h0;  // 32'h100bc775;
    ram_cell[     188] = 32'h0;  // 32'h11c60095;
    ram_cell[     189] = 32'h0;  // 32'h0c3c0e91;
    ram_cell[     190] = 32'h0;  // 32'h73b25d72;
    ram_cell[     191] = 32'h0;  // 32'hff577268;
    ram_cell[     192] = 32'h0;  // 32'h84ac2a7f;
    ram_cell[     193] = 32'h0;  // 32'hc3017f9c;
    ram_cell[     194] = 32'h0;  // 32'h85031707;
    ram_cell[     195] = 32'h0;  // 32'hde04cc52;
    ram_cell[     196] = 32'h0;  // 32'h12c0070e;
    ram_cell[     197] = 32'h0;  // 32'hda1442b1;
    ram_cell[     198] = 32'h0;  // 32'hc661084c;
    ram_cell[     199] = 32'h0;  // 32'h43384c20;
    ram_cell[     200] = 32'h0;  // 32'hd831ab58;
    ram_cell[     201] = 32'h0;  // 32'h58a09163;
    ram_cell[     202] = 32'h0;  // 32'h4c050837;
    ram_cell[     203] = 32'h0;  // 32'h21f65ecb;
    ram_cell[     204] = 32'h0;  // 32'h9624de07;
    ram_cell[     205] = 32'h0;  // 32'h15cf4d66;
    ram_cell[     206] = 32'h0;  // 32'h5dad15fd;
    ram_cell[     207] = 32'h0;  // 32'h14b728b3;
    ram_cell[     208] = 32'h0;  // 32'h43f714da;
    ram_cell[     209] = 32'h0;  // 32'h4b39d52f;
    ram_cell[     210] = 32'h0;  // 32'he7b7f29d;
    ram_cell[     211] = 32'h0;  // 32'h54f69c4e;
    ram_cell[     212] = 32'h0;  // 32'h1e613e19;
    ram_cell[     213] = 32'h0;  // 32'h85bfe765;
    ram_cell[     214] = 32'h0;  // 32'h0c0e8718;
    ram_cell[     215] = 32'h0;  // 32'h7e976f83;
    ram_cell[     216] = 32'h0;  // 32'h7cd75f86;
    ram_cell[     217] = 32'h0;  // 32'hea75af0b;
    ram_cell[     218] = 32'h0;  // 32'h8a37bf5a;
    ram_cell[     219] = 32'h0;  // 32'hd2100bd8;
    ram_cell[     220] = 32'h0;  // 32'haa5e7252;
    ram_cell[     221] = 32'h0;  // 32'h6b5b673a;
    ram_cell[     222] = 32'h0;  // 32'h6f0741f4;
    ram_cell[     223] = 32'h0;  // 32'hc8c26a1a;
    ram_cell[     224] = 32'h0;  // 32'h650e6515;
    ram_cell[     225] = 32'h0;  // 32'h23bfadce;
    ram_cell[     226] = 32'h0;  // 32'hea2d0fe7;
    ram_cell[     227] = 32'h0;  // 32'h55ef72ea;
    ram_cell[     228] = 32'h0;  // 32'h747a74f2;
    ram_cell[     229] = 32'h0;  // 32'hc352286e;
    ram_cell[     230] = 32'h0;  // 32'hfae23a81;
    ram_cell[     231] = 32'h0;  // 32'h8b0c42ee;
    ram_cell[     232] = 32'h0;  // 32'h6461ae4c;
    ram_cell[     233] = 32'h0;  // 32'hf28e6780;
    ram_cell[     234] = 32'h0;  // 32'hde1c1bef;
    ram_cell[     235] = 32'h0;  // 32'hbcc3dda8;
    ram_cell[     236] = 32'h0;  // 32'hecaa50ee;
    ram_cell[     237] = 32'h0;  // 32'hf0bbe8dd;
    ram_cell[     238] = 32'h0;  // 32'hd3e36921;
    ram_cell[     239] = 32'h0;  // 32'h88709362;
    ram_cell[     240] = 32'h0;  // 32'h8f0e7b8f;
    ram_cell[     241] = 32'h0;  // 32'hbce11d3e;
    ram_cell[     242] = 32'h0;  // 32'h63aa922a;
    ram_cell[     243] = 32'h0;  // 32'hf51d9747;
    ram_cell[     244] = 32'h0;  // 32'h04c4d07a;
    ram_cell[     245] = 32'h0;  // 32'h075cdf3f;
    ram_cell[     246] = 32'h0;  // 32'hec034846;
    ram_cell[     247] = 32'h0;  // 32'h9e6046f2;
    ram_cell[     248] = 32'h0;  // 32'h563650c2;
    ram_cell[     249] = 32'h0;  // 32'h8a212c7a;
    ram_cell[     250] = 32'h0;  // 32'hb05a3ff6;
    ram_cell[     251] = 32'h0;  // 32'h66911a73;
    ram_cell[     252] = 32'h0;  // 32'hee0b2e31;
    ram_cell[     253] = 32'h0;  // 32'h65e62856;
    ram_cell[     254] = 32'h0;  // 32'h64380c48;
    ram_cell[     255] = 32'h0;  // 32'hb38965eb;
    // src matrix A
    ram_cell[     256] = 32'hcdb99e1d;
    ram_cell[     257] = 32'h3630b58a;
    ram_cell[     258] = 32'hb1df2d11;
    ram_cell[     259] = 32'hdac93b03;
    ram_cell[     260] = 32'hcbbfd78d;
    ram_cell[     261] = 32'h3b11116c;
    ram_cell[     262] = 32'h171f7680;
    ram_cell[     263] = 32'hd6d623c5;
    ram_cell[     264] = 32'hfda338da;
    ram_cell[     265] = 32'h2ed044a8;
    ram_cell[     266] = 32'hbfc63cb1;
    ram_cell[     267] = 32'h1fd0f92f;
    ram_cell[     268] = 32'h4372b921;
    ram_cell[     269] = 32'hc9f40af0;
    ram_cell[     270] = 32'hb8e90bdc;
    ram_cell[     271] = 32'h5f470816;
    ram_cell[     272] = 32'h6bbd9e90;
    ram_cell[     273] = 32'h1d66206d;
    ram_cell[     274] = 32'hf688e177;
    ram_cell[     275] = 32'h30af8905;
    ram_cell[     276] = 32'hca03e7b5;
    ram_cell[     277] = 32'he1412b80;
    ram_cell[     278] = 32'h6593f949;
    ram_cell[     279] = 32'h50b78ce5;
    ram_cell[     280] = 32'h342f5024;
    ram_cell[     281] = 32'h70a36be9;
    ram_cell[     282] = 32'ha8b93264;
    ram_cell[     283] = 32'h202bc5ed;
    ram_cell[     284] = 32'hafc7aec1;
    ram_cell[     285] = 32'h969a1dc1;
    ram_cell[     286] = 32'h587fb538;
    ram_cell[     287] = 32'h0d6b7382;
    ram_cell[     288] = 32'heb28ea44;
    ram_cell[     289] = 32'h636b6279;
    ram_cell[     290] = 32'h8eb95d64;
    ram_cell[     291] = 32'h53f15b14;
    ram_cell[     292] = 32'he0b0eded;
    ram_cell[     293] = 32'h841da49b;
    ram_cell[     294] = 32'h057ccaa3;
    ram_cell[     295] = 32'h92ba76cb;
    ram_cell[     296] = 32'h24ff7721;
    ram_cell[     297] = 32'h7b75ca02;
    ram_cell[     298] = 32'hfad3af70;
    ram_cell[     299] = 32'h9023d8dd;
    ram_cell[     300] = 32'h4c3defe7;
    ram_cell[     301] = 32'h861c9ebf;
    ram_cell[     302] = 32'ha929a4ed;
    ram_cell[     303] = 32'hd31c59b9;
    ram_cell[     304] = 32'hc45969a3;
    ram_cell[     305] = 32'h300ca050;
    ram_cell[     306] = 32'h7cdd28c8;
    ram_cell[     307] = 32'hde03a12f;
    ram_cell[     308] = 32'he882b85d;
    ram_cell[     309] = 32'h94b130e9;
    ram_cell[     310] = 32'hebfb24af;
    ram_cell[     311] = 32'h839edb32;
    ram_cell[     312] = 32'hda87e320;
    ram_cell[     313] = 32'hd2190079;
    ram_cell[     314] = 32'h4e856319;
    ram_cell[     315] = 32'h3fe6755b;
    ram_cell[     316] = 32'ha0c6ab5b;
    ram_cell[     317] = 32'h4ff0ee10;
    ram_cell[     318] = 32'ha7f20cf4;
    ram_cell[     319] = 32'h3d43ab29;
    ram_cell[     320] = 32'hd1e11263;
    ram_cell[     321] = 32'h9b805709;
    ram_cell[     322] = 32'h6af15373;
    ram_cell[     323] = 32'h8f9fd7c4;
    ram_cell[     324] = 32'h76dcf0fd;
    ram_cell[     325] = 32'h43050eda;
    ram_cell[     326] = 32'h1e5c6c55;
    ram_cell[     327] = 32'he859d24b;
    ram_cell[     328] = 32'hb33d2f2b;
    ram_cell[     329] = 32'h9cb29f46;
    ram_cell[     330] = 32'hc5cce0a1;
    ram_cell[     331] = 32'h8b47db9c;
    ram_cell[     332] = 32'hd54de4d5;
    ram_cell[     333] = 32'he462fe33;
    ram_cell[     334] = 32'hde002559;
    ram_cell[     335] = 32'h84d36b83;
    ram_cell[     336] = 32'h0ecc25b2;
    ram_cell[     337] = 32'hbb6fcbff;
    ram_cell[     338] = 32'h7a8f27de;
    ram_cell[     339] = 32'ha1cfff6f;
    ram_cell[     340] = 32'h93d941f4;
    ram_cell[     341] = 32'h76646e5f;
    ram_cell[     342] = 32'h6ab10cf7;
    ram_cell[     343] = 32'h2a752509;
    ram_cell[     344] = 32'hca6f03b2;
    ram_cell[     345] = 32'h3471531f;
    ram_cell[     346] = 32'hb0cb0b4b;
    ram_cell[     347] = 32'h6df2f7c7;
    ram_cell[     348] = 32'h5f8cfef3;
    ram_cell[     349] = 32'hfe47cd90;
    ram_cell[     350] = 32'h27cf78d5;
    ram_cell[     351] = 32'h62fe4832;
    ram_cell[     352] = 32'h912e8f57;
    ram_cell[     353] = 32'hc55b6e88;
    ram_cell[     354] = 32'h36acd172;
    ram_cell[     355] = 32'heaa0b364;
    ram_cell[     356] = 32'h6ff51293;
    ram_cell[     357] = 32'he023448c;
    ram_cell[     358] = 32'h27db4332;
    ram_cell[     359] = 32'h9d861b4e;
    ram_cell[     360] = 32'h513642f6;
    ram_cell[     361] = 32'h0313e80a;
    ram_cell[     362] = 32'ha0174631;
    ram_cell[     363] = 32'h20c7baa5;
    ram_cell[     364] = 32'hce4720d2;
    ram_cell[     365] = 32'h7cd93cdf;
    ram_cell[     366] = 32'hb7a20784;
    ram_cell[     367] = 32'h03074455;
    ram_cell[     368] = 32'h09d78a86;
    ram_cell[     369] = 32'h55918b37;
    ram_cell[     370] = 32'h10578102;
    ram_cell[     371] = 32'h57db0750;
    ram_cell[     372] = 32'h64eaab49;
    ram_cell[     373] = 32'h79c2ec55;
    ram_cell[     374] = 32'h96d9a81b;
    ram_cell[     375] = 32'h9b9d1db3;
    ram_cell[     376] = 32'ha1c90aa4;
    ram_cell[     377] = 32'h556f9ab2;
    ram_cell[     378] = 32'h18b94761;
    ram_cell[     379] = 32'hf8e7fd78;
    ram_cell[     380] = 32'h8d0c0409;
    ram_cell[     381] = 32'h05ae4b58;
    ram_cell[     382] = 32'h3e40f2e6;
    ram_cell[     383] = 32'h2b14717a;
    ram_cell[     384] = 32'h88f406a0;
    ram_cell[     385] = 32'h1e75ede9;
    ram_cell[     386] = 32'h149a608c;
    ram_cell[     387] = 32'he5d9d77d;
    ram_cell[     388] = 32'haeaced25;
    ram_cell[     389] = 32'hf45f1e10;
    ram_cell[     390] = 32'hd8f2ead5;
    ram_cell[     391] = 32'h317fdfd5;
    ram_cell[     392] = 32'ha8ca01b2;
    ram_cell[     393] = 32'h003812f6;
    ram_cell[     394] = 32'h73b0c87b;
    ram_cell[     395] = 32'hc5ea0d6d;
    ram_cell[     396] = 32'hab353b20;
    ram_cell[     397] = 32'h6280a446;
    ram_cell[     398] = 32'h36648837;
    ram_cell[     399] = 32'h21dd184f;
    ram_cell[     400] = 32'he8f803ca;
    ram_cell[     401] = 32'he45d9e1f;
    ram_cell[     402] = 32'h00be1f85;
    ram_cell[     403] = 32'h1703b29d;
    ram_cell[     404] = 32'hf2e7fe1c;
    ram_cell[     405] = 32'he555cf44;
    ram_cell[     406] = 32'h2ca1e1c0;
    ram_cell[     407] = 32'hcc748d44;
    ram_cell[     408] = 32'h84c2979c;
    ram_cell[     409] = 32'h8baca171;
    ram_cell[     410] = 32'hdead8845;
    ram_cell[     411] = 32'h62d27efe;
    ram_cell[     412] = 32'h7c02dee4;
    ram_cell[     413] = 32'h27000107;
    ram_cell[     414] = 32'h1ba27e36;
    ram_cell[     415] = 32'h5793e933;
    ram_cell[     416] = 32'had165e81;
    ram_cell[     417] = 32'h4a5b3619;
    ram_cell[     418] = 32'h1d89b114;
    ram_cell[     419] = 32'hd6dd9784;
    ram_cell[     420] = 32'h581a0af4;
    ram_cell[     421] = 32'h7f4ddc36;
    ram_cell[     422] = 32'haefeec6e;
    ram_cell[     423] = 32'h649f8603;
    ram_cell[     424] = 32'h72c2520d;
    ram_cell[     425] = 32'h22b12f3c;
    ram_cell[     426] = 32'hf57083fe;
    ram_cell[     427] = 32'hed35a1c3;
    ram_cell[     428] = 32'h063f2907;
    ram_cell[     429] = 32'hb44f5314;
    ram_cell[     430] = 32'h9937cc21;
    ram_cell[     431] = 32'h92a34997;
    ram_cell[     432] = 32'haffaf0de;
    ram_cell[     433] = 32'hb618f92f;
    ram_cell[     434] = 32'h601d0cad;
    ram_cell[     435] = 32'hc0b8acfe;
    ram_cell[     436] = 32'h80b98ce6;
    ram_cell[     437] = 32'h988587d1;
    ram_cell[     438] = 32'h90b9d7b7;
    ram_cell[     439] = 32'hc39c2206;
    ram_cell[     440] = 32'ha0add570;
    ram_cell[     441] = 32'ha3492d35;
    ram_cell[     442] = 32'h6ea50ffa;
    ram_cell[     443] = 32'h0984c70b;
    ram_cell[     444] = 32'hdac3815c;
    ram_cell[     445] = 32'h9e91abcb;
    ram_cell[     446] = 32'he220a546;
    ram_cell[     447] = 32'h60be20ba;
    ram_cell[     448] = 32'h72ff0828;
    ram_cell[     449] = 32'hbba77f2d;
    ram_cell[     450] = 32'h9504dcd9;
    ram_cell[     451] = 32'h5015b821;
    ram_cell[     452] = 32'hecefed56;
    ram_cell[     453] = 32'hf5cc83b6;
    ram_cell[     454] = 32'hc0449c89;
    ram_cell[     455] = 32'h4c94af39;
    ram_cell[     456] = 32'hcb2d458a;
    ram_cell[     457] = 32'hd943db18;
    ram_cell[     458] = 32'hd247e83e;
    ram_cell[     459] = 32'h11db1016;
    ram_cell[     460] = 32'h10de3fea;
    ram_cell[     461] = 32'hb0f3e7c6;
    ram_cell[     462] = 32'hb73c06a0;
    ram_cell[     463] = 32'h686ec8f4;
    ram_cell[     464] = 32'h29f755ab;
    ram_cell[     465] = 32'h5198673a;
    ram_cell[     466] = 32'he0ef10bf;
    ram_cell[     467] = 32'ha72be0dc;
    ram_cell[     468] = 32'hf0e67362;
    ram_cell[     469] = 32'h4aa8cc11;
    ram_cell[     470] = 32'hf744e2f7;
    ram_cell[     471] = 32'hff5a962a;
    ram_cell[     472] = 32'h51921e36;
    ram_cell[     473] = 32'he287cd92;
    ram_cell[     474] = 32'h10bdaf56;
    ram_cell[     475] = 32'h667d0267;
    ram_cell[     476] = 32'h10a907c3;
    ram_cell[     477] = 32'h599a2ddf;
    ram_cell[     478] = 32'hd809ef40;
    ram_cell[     479] = 32'hf39c6e6f;
    ram_cell[     480] = 32'hc62770ca;
    ram_cell[     481] = 32'h2c834816;
    ram_cell[     482] = 32'hdc05114b;
    ram_cell[     483] = 32'heeeb2ca7;
    ram_cell[     484] = 32'hba07414c;
    ram_cell[     485] = 32'h37006096;
    ram_cell[     486] = 32'h23549715;
    ram_cell[     487] = 32'haa8317b4;
    ram_cell[     488] = 32'h107222e7;
    ram_cell[     489] = 32'h8212b80f;
    ram_cell[     490] = 32'h8a934bcb;
    ram_cell[     491] = 32'h30d2d769;
    ram_cell[     492] = 32'h98ff395b;
    ram_cell[     493] = 32'h1de339bf;
    ram_cell[     494] = 32'h784e2de5;
    ram_cell[     495] = 32'h45424a94;
    ram_cell[     496] = 32'hca5758f8;
    ram_cell[     497] = 32'h779747db;
    ram_cell[     498] = 32'h8722462c;
    ram_cell[     499] = 32'h6d3c9128;
    ram_cell[     500] = 32'h9da25bfb;
    ram_cell[     501] = 32'h54bf93fd;
    ram_cell[     502] = 32'h7d5fbe9b;
    ram_cell[     503] = 32'h2722f8c1;
    ram_cell[     504] = 32'h792f5b4e;
    ram_cell[     505] = 32'h4ee82df9;
    ram_cell[     506] = 32'h2234a61d;
    ram_cell[     507] = 32'h88a20af8;
    ram_cell[     508] = 32'h2f9174fc;
    ram_cell[     509] = 32'h9b55207e;
    ram_cell[     510] = 32'h50bfb44d;
    ram_cell[     511] = 32'h284fca37;
    // src matrix B
    ram_cell[     512] = 32'h21a06f1f;
    ram_cell[     513] = 32'h9173de4e;
    ram_cell[     514] = 32'h3794ca6f;
    ram_cell[     515] = 32'h68dd1d93;
    ram_cell[     516] = 32'hc8047a6b;
    ram_cell[     517] = 32'ha34056b2;
    ram_cell[     518] = 32'h541f18f2;
    ram_cell[     519] = 32'hd1a18d2e;
    ram_cell[     520] = 32'h538181b5;
    ram_cell[     521] = 32'h96366cc6;
    ram_cell[     522] = 32'h8ef04a75;
    ram_cell[     523] = 32'h005e4ca5;
    ram_cell[     524] = 32'h7c656870;
    ram_cell[     525] = 32'he6ed2ff6;
    ram_cell[     526] = 32'h43c4ff67;
    ram_cell[     527] = 32'h8455b5bf;
    ram_cell[     528] = 32'h9ce62328;
    ram_cell[     529] = 32'h0728d273;
    ram_cell[     530] = 32'h87da9967;
    ram_cell[     531] = 32'h9d1126aa;
    ram_cell[     532] = 32'hb18749d7;
    ram_cell[     533] = 32'hae36b03a;
    ram_cell[     534] = 32'hc5f1b864;
    ram_cell[     535] = 32'hc2df7315;
    ram_cell[     536] = 32'h67a4bb2f;
    ram_cell[     537] = 32'h38f62f93;
    ram_cell[     538] = 32'hdf5efeb7;
    ram_cell[     539] = 32'h28694b71;
    ram_cell[     540] = 32'hf2fb85cc;
    ram_cell[     541] = 32'hbd21d351;
    ram_cell[     542] = 32'h45f355fa;
    ram_cell[     543] = 32'h13a3fede;
    ram_cell[     544] = 32'h9a89a761;
    ram_cell[     545] = 32'h76b40287;
    ram_cell[     546] = 32'h53f97129;
    ram_cell[     547] = 32'h4e865e8c;
    ram_cell[     548] = 32'h33366630;
    ram_cell[     549] = 32'hc4f91df9;
    ram_cell[     550] = 32'h04b31698;
    ram_cell[     551] = 32'hfe823a16;
    ram_cell[     552] = 32'heeece094;
    ram_cell[     553] = 32'hcce814d9;
    ram_cell[     554] = 32'hed71438a;
    ram_cell[     555] = 32'h0f01d5a9;
    ram_cell[     556] = 32'h6f3bf5bd;
    ram_cell[     557] = 32'h167e9924;
    ram_cell[     558] = 32'hb428d867;
    ram_cell[     559] = 32'h0d1e7d56;
    ram_cell[     560] = 32'h184c620e;
    ram_cell[     561] = 32'haa98b23f;
    ram_cell[     562] = 32'h95a8f6ef;
    ram_cell[     563] = 32'h4ab3161c;
    ram_cell[     564] = 32'hd33da2d9;
    ram_cell[     565] = 32'h4090cf49;
    ram_cell[     566] = 32'hfa5f2f09;
    ram_cell[     567] = 32'h298fc302;
    ram_cell[     568] = 32'hda53665a;
    ram_cell[     569] = 32'h6ff2bb67;
    ram_cell[     570] = 32'h90d38d3e;
    ram_cell[     571] = 32'h447e1771;
    ram_cell[     572] = 32'hcd7bf27a;
    ram_cell[     573] = 32'hc5d869b1;
    ram_cell[     574] = 32'h98048e79;
    ram_cell[     575] = 32'h72ab12e2;
    ram_cell[     576] = 32'hd2501d2a;
    ram_cell[     577] = 32'he03cc77c;
    ram_cell[     578] = 32'h7712f183;
    ram_cell[     579] = 32'h724f8297;
    ram_cell[     580] = 32'hc4f50d87;
    ram_cell[     581] = 32'hd5826d81;
    ram_cell[     582] = 32'hf4755f53;
    ram_cell[     583] = 32'h72947238;
    ram_cell[     584] = 32'hd70a7fda;
    ram_cell[     585] = 32'h851022b4;
    ram_cell[     586] = 32'h0c96dc96;
    ram_cell[     587] = 32'h9e3ff063;
    ram_cell[     588] = 32'h8a8c27be;
    ram_cell[     589] = 32'h6007b09b;
    ram_cell[     590] = 32'ha81423e9;
    ram_cell[     591] = 32'h1953224f;
    ram_cell[     592] = 32'h9924ff2f;
    ram_cell[     593] = 32'hc8781d3b;
    ram_cell[     594] = 32'h001257f9;
    ram_cell[     595] = 32'hbc4ecb48;
    ram_cell[     596] = 32'hd890a957;
    ram_cell[     597] = 32'hfb896f64;
    ram_cell[     598] = 32'he51c9a96;
    ram_cell[     599] = 32'h444ece3e;
    ram_cell[     600] = 32'h0ba9bbc3;
    ram_cell[     601] = 32'h426eeba1;
    ram_cell[     602] = 32'h4ce809f6;
    ram_cell[     603] = 32'h246afdf7;
    ram_cell[     604] = 32'h9066f84b;
    ram_cell[     605] = 32'h2012488a;
    ram_cell[     606] = 32'h761da6de;
    ram_cell[     607] = 32'h08d83766;
    ram_cell[     608] = 32'h9fe685ec;
    ram_cell[     609] = 32'h44543586;
    ram_cell[     610] = 32'h8b595aac;
    ram_cell[     611] = 32'h7ed0e7c1;
    ram_cell[     612] = 32'h975aaddf;
    ram_cell[     613] = 32'h810bae52;
    ram_cell[     614] = 32'hac129dc5;
    ram_cell[     615] = 32'h723c5554;
    ram_cell[     616] = 32'hecbca52a;
    ram_cell[     617] = 32'h6aeffa08;
    ram_cell[     618] = 32'h1c1a5bf9;
    ram_cell[     619] = 32'hfd4cb00b;
    ram_cell[     620] = 32'ha0e118f3;
    ram_cell[     621] = 32'hade9ad25;
    ram_cell[     622] = 32'hc263b129;
    ram_cell[     623] = 32'heb069043;
    ram_cell[     624] = 32'hdc7690e2;
    ram_cell[     625] = 32'h2d245ae5;
    ram_cell[     626] = 32'h3a1fdb0a;
    ram_cell[     627] = 32'h5c739b99;
    ram_cell[     628] = 32'h3c5d06fd;
    ram_cell[     629] = 32'h355470fd;
    ram_cell[     630] = 32'h1ad1ad08;
    ram_cell[     631] = 32'h17579807;
    ram_cell[     632] = 32'haa7e1519;
    ram_cell[     633] = 32'h8bec5ce2;
    ram_cell[     634] = 32'h3747cdcb;
    ram_cell[     635] = 32'hbefda70b;
    ram_cell[     636] = 32'h0ee06917;
    ram_cell[     637] = 32'hfcb37669;
    ram_cell[     638] = 32'h79021bf0;
    ram_cell[     639] = 32'hc699873c;
    ram_cell[     640] = 32'h599c3ead;
    ram_cell[     641] = 32'h04cacf2e;
    ram_cell[     642] = 32'h96362088;
    ram_cell[     643] = 32'h52577669;
    ram_cell[     644] = 32'hd6b80587;
    ram_cell[     645] = 32'h40451499;
    ram_cell[     646] = 32'he0acc3e6;
    ram_cell[     647] = 32'h0f8f91a5;
    ram_cell[     648] = 32'h6c3963a1;
    ram_cell[     649] = 32'h908b4ba9;
    ram_cell[     650] = 32'h7cdc7959;
    ram_cell[     651] = 32'h1868ad35;
    ram_cell[     652] = 32'h210ce773;
    ram_cell[     653] = 32'h4159799e;
    ram_cell[     654] = 32'h1ed2d9a3;
    ram_cell[     655] = 32'h87293014;
    ram_cell[     656] = 32'he14b9e82;
    ram_cell[     657] = 32'h48150ded;
    ram_cell[     658] = 32'h369e186b;
    ram_cell[     659] = 32'hedc9c15d;
    ram_cell[     660] = 32'h3a2c9b36;
    ram_cell[     661] = 32'h150c07ed;
    ram_cell[     662] = 32'hc286061e;
    ram_cell[     663] = 32'h8d7f87ba;
    ram_cell[     664] = 32'h58818d37;
    ram_cell[     665] = 32'hb3bd871f;
    ram_cell[     666] = 32'h6ecffb03;
    ram_cell[     667] = 32'h4f42bb12;
    ram_cell[     668] = 32'h516cb499;
    ram_cell[     669] = 32'h592fd33c;
    ram_cell[     670] = 32'h867f6c39;
    ram_cell[     671] = 32'h129162d8;
    ram_cell[     672] = 32'hc8a33544;
    ram_cell[     673] = 32'h4a7c00ca;
    ram_cell[     674] = 32'h0b1757d0;
    ram_cell[     675] = 32'hb16b38c8;
    ram_cell[     676] = 32'hdb607eda;
    ram_cell[     677] = 32'h65fa3cb7;
    ram_cell[     678] = 32'h822d131a;
    ram_cell[     679] = 32'h4240fbfa;
    ram_cell[     680] = 32'heaea04ca;
    ram_cell[     681] = 32'hf1985353;
    ram_cell[     682] = 32'h24d7a5fb;
    ram_cell[     683] = 32'h76b661b3;
    ram_cell[     684] = 32'h6d8ce2c0;
    ram_cell[     685] = 32'hef3f785f;
    ram_cell[     686] = 32'ha5d5f58f;
    ram_cell[     687] = 32'h40bb7a3f;
    ram_cell[     688] = 32'h5b51bda6;
    ram_cell[     689] = 32'h0a201f64;
    ram_cell[     690] = 32'h7dbdd0a9;
    ram_cell[     691] = 32'hca0f5d67;
    ram_cell[     692] = 32'hc79f8046;
    ram_cell[     693] = 32'h545c2d5e;
    ram_cell[     694] = 32'h01fad0e2;
    ram_cell[     695] = 32'h0f3dcd69;
    ram_cell[     696] = 32'hf493c14f;
    ram_cell[     697] = 32'h25b78476;
    ram_cell[     698] = 32'hb67e227b;
    ram_cell[     699] = 32'h259e860a;
    ram_cell[     700] = 32'hf00a8f50;
    ram_cell[     701] = 32'h3940cd4b;
    ram_cell[     702] = 32'h3ac96b04;
    ram_cell[     703] = 32'h96584982;
    ram_cell[     704] = 32'h332c8fad;
    ram_cell[     705] = 32'h620b4599;
    ram_cell[     706] = 32'h947c35de;
    ram_cell[     707] = 32'hb7e39be4;
    ram_cell[     708] = 32'h6a291ee1;
    ram_cell[     709] = 32'hbec313a2;
    ram_cell[     710] = 32'hfab31094;
    ram_cell[     711] = 32'h5f14ac50;
    ram_cell[     712] = 32'h36d78612;
    ram_cell[     713] = 32'h68d8b2a1;
    ram_cell[     714] = 32'hed3c7ab7;
    ram_cell[     715] = 32'h53f77e3b;
    ram_cell[     716] = 32'h13fd7e6f;
    ram_cell[     717] = 32'h7395b275;
    ram_cell[     718] = 32'hf93da437;
    ram_cell[     719] = 32'h6b1b4c87;
    ram_cell[     720] = 32'h4ad7375d;
    ram_cell[     721] = 32'h7cc0676b;
    ram_cell[     722] = 32'h934d9a04;
    ram_cell[     723] = 32'h4ca69d0d;
    ram_cell[     724] = 32'hd5544f71;
    ram_cell[     725] = 32'hd7a85a79;
    ram_cell[     726] = 32'h3f5a9cc4;
    ram_cell[     727] = 32'hde5970ff;
    ram_cell[     728] = 32'h6c34d47d;
    ram_cell[     729] = 32'h55a59d40;
    ram_cell[     730] = 32'h4166d79f;
    ram_cell[     731] = 32'h3e0f4085;
    ram_cell[     732] = 32'h1eceab55;
    ram_cell[     733] = 32'ha2cc7700;
    ram_cell[     734] = 32'hf2fc04df;
    ram_cell[     735] = 32'h2e191769;
    ram_cell[     736] = 32'h4917317f;
    ram_cell[     737] = 32'hf3da8db3;
    ram_cell[     738] = 32'h7b93dd93;
    ram_cell[     739] = 32'h3288d0f1;
    ram_cell[     740] = 32'h0842ba37;
    ram_cell[     741] = 32'hecb682b2;
    ram_cell[     742] = 32'h096b10e9;
    ram_cell[     743] = 32'h734670b3;
    ram_cell[     744] = 32'h34e5987a;
    ram_cell[     745] = 32'h487fe1d2;
    ram_cell[     746] = 32'h0257d696;
    ram_cell[     747] = 32'h1982374b;
    ram_cell[     748] = 32'h847c8712;
    ram_cell[     749] = 32'h52a018ca;
    ram_cell[     750] = 32'h3c33876b;
    ram_cell[     751] = 32'h72e0fc8e;
    ram_cell[     752] = 32'h302dd0a3;
    ram_cell[     753] = 32'h416dc621;
    ram_cell[     754] = 32'hcd204d61;
    ram_cell[     755] = 32'ha5b2404a;
    ram_cell[     756] = 32'h66856300;
    ram_cell[     757] = 32'h2f49fed7;
    ram_cell[     758] = 32'h0beeaf67;
    ram_cell[     759] = 32'hcd0ce225;
    ram_cell[     760] = 32'h28209488;
    ram_cell[     761] = 32'hc84bbe6c;
    ram_cell[     762] = 32'h2424a3fb;
    ram_cell[     763] = 32'hc23c2bec;
    ram_cell[     764] = 32'hd652eaa3;
    ram_cell[     765] = 32'hb80adfc5;
    ram_cell[     766] = 32'hc460a399;
    ram_cell[     767] = 32'h785940da;
end

endmodule

